`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   17:34:19 09/11/2015
// Design Name:   Lab9_1
// Module Name:   G:/HP LAB/file/Lab9_1/Lab9_1_test.v
// Project Name:  Lab9_1
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Lab9_1
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module Lab9_1_test;

	// Inputs
	reg clk;
	reg reset;
	reg [15:0] audio_in_left;
	reg [15:0] audio_in_right;

	// Outputs
	wire audio_appsel;
	wire audio_sysclk;
	wire audio_bck;
	wire audio_ws;
	wire audio_data;

	// Instantiate the Unit Under Test (UUT)
	Lab9_1 uut (
		.clk(clk), 
		.reset(reset), 
		.audio_in_left(audio_in_left), 
		.audio_in_right(audio_in_right), 
		.audio_appsel(audio_appsel), 
		.audio_sysclk(audio_sysclk), 
		.audio_bck(audio_bck), 
		.audio_ws(audio_ws), 
		.audio_data(audio_data)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 0;
		audio_in_left = 16'h3FFF;
		audio_in_right = 16'hC000;

		// Wait 100 ns for global reset to finish
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;reset = 1;  //100 
		// Add stimulus here
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000

#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
		
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//100
		#25 clk =1;
		#25 clk =0;
      #25 clk =1;
		#25 clk =0;//1000
	end
      
endmodule

